// this file is placeholder for common code
